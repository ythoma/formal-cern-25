library ieee;
use ieee.std_logic_1164.all;

entity psl_sequence is
    generic (
        EXPECT_FAIL : boolean := false
    );
    port (
        clk : in std_logic
    );
end entity psl_sequence;

architecture psl of psl_sequence is

    signal a, b: std_logic;

begin

    -- All is sensitive to rising edge of clk
    default clock is rising_edge(clk);


    --                                          012345678901
    seq_a : entity work.sequencer generic map ("-____-__-___") port map (clk, a);
    seq_b : entity work.sequencer generic map ("__-__-___-__") port map (clk, b);

    assert_success1a: assert (a -> not b);
    assert_success1b: assert (b -> not a);
 
    gen_fail : if EXPECT_FAIL generate
        assert_fail1: assert not(a and b);
        assert_fail2: assert always not(a and b);
        assert_fail3: assert never (a and b);
    end generate;

end architecture psl;
