library ieee;

package bpm_pkg is

    constant CONST_MIN_DT_TIME           : integer := 4;
    constant CONST_MIN_OT_TIME           : integer := 4;

end package;